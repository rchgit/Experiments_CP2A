`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:58:32 01/29/2014 
// Design Name: 
// Module Name:    DRAP_REGFILE 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//parameterized register File
module DRAP_REGFILE
#(
parameter B = 32, //number of bits
W = 5 //number of address bits
)
(input wire clk,
input wire rst, wr_en,
input wire [W-1:0] r_addr1, r_addr2, w_addr,
input wire [B-1:0] w_data,
output wire [B-1:0] r_data1, r_data2);
reg [B-1:0] array_reg [2**W-1:0];// = 32'b00000000_00000000_00000000_00000000;
always @(posedge clk, posedge rst)
	if (rst)
		begin
			array_reg[5'b00000] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00001] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00010] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00011] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00100] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00101] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00110] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b00111] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01000] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01001] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01010] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01011] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01100] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01101] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01110] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b01111] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10000] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10001] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10010] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10011] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10100] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10101] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10110] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b10111] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11000] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11001] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11010] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11011] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11100] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11101] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11110] <= 32'b00000000_00000000_00000000_00000000;
			array_reg[5'b11111] <= 32'b00000000_00000000_00000000_00000000;
		end
	else
		if (wr_en)
			array_reg[w_addr] <=w_data;
// read operation
assign r_data1 = array_reg[r_addr1];
assign r_data2 = array_reg[r_addr2];
endmodule
